15 gid=1161177
15 uid=1161177
30 mtime=1483662701.000000001
20 ctime=1483662701
20 atime=1483662701
