15 gid=1161177
15 uid=1161177
30 mtime=1482221023.000000001
20 ctime=1482221023
20 atime=1482221023
