15 gid=1161177
15 uid=1161177
30 mtime=1485439165.000000001
20 ctime=1485439165
20 atime=1485439165
