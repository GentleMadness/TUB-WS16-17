15 gid=1161177
15 uid=1161177
30 mtime=1483667645.000000001
20 ctime=1483667645
20 atime=1483667645
