15 gid=1161177
15 uid=1161177
30 mtime=1484929677.000000001
20 ctime=1484929677
20 atime=1484929677
