15 gid=1161177
15 uid=1161177
30 mtime=1484831206.000000001
20 ctime=1484831206
20 atime=1484831206
