15 gid=1161177
15 uid=1161177
30 mtime=1485441620.000000001
20 ctime=1485441620
20 atime=1485441620
