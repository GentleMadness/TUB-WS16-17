15 gid=1161177
15 uid=1161177
30 mtime=1484939937.000000001
20 ctime=1484939937
20 atime=1484939937
