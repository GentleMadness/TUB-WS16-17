15 gid=1161177
15 uid=1161177
30 mtime=1482220738.000000001
20 ctime=1482220738
20 atime=1482220738
