15 gid=1161177
15 uid=1161177
30 mtime=1482220840.000000001
20 ctime=1482220840
20 atime=1482220840
