15 gid=1161177
15 uid=1161177
30 mtime=1485382555.000000001
20 ctime=1485382555
20 atime=1485382555
