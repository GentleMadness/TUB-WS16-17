15 gid=1161177
15 uid=1161177
30 mtime=1483668090.000000001
20 ctime=1483668090
20 atime=1483668090
